402
411
#
#

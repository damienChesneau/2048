401
433
#
#
